magic
tech scmos
timestamp 1701770819
<< polysilicon >>
rect 143 962 511 964
rect 143 181 145 962
rect 265 605 323 607
rect 265 245 267 605
rect 145 107 255 109
rect 142 -1157 144 35
rect 253 -186 255 107
rect 253 -188 322 -186
rect 435 -1061 542 -1059
rect 142 -1159 336 -1157
rect 435 -1203 437 -1061
rect 445 -1131 542 -1129
rect 445 -1275 447 -1131
rect 439 -1277 447 -1275
rect 466 -1203 542 -1201
rect 466 -1346 468 -1203
rect 439 -1348 468 -1346
rect 501 -1274 542 -1272
rect 501 -1417 503 -1274
rect 438 -1419 503 -1417
<< polycontact >>
rect 511 960 515 964
rect 323 604 327 608
rect 264 241 268 245
rect 142 177 146 181
rect 141 106 145 110
rect 141 35 145 39
rect 322 -189 326 -185
rect 336 -1160 340 -1156
rect 542 -1062 546 -1058
rect 434 -1207 438 -1203
rect 435 -1278 439 -1274
rect 542 -1133 546 -1129
rect 435 -1349 439 -1345
rect 542 -1204 546 -1200
rect 434 -1420 438 -1416
rect 542 -1275 546 -1271
<< metal1 >>
rect 515 960 516 964
rect 440 952 521 956
rect -553 857 335 861
rect 440 860 444 952
rect -553 -145 -549 857
rect 416 856 444 860
rect -493 786 335 790
rect -493 -100 -489 786
rect 418 785 508 789
rect 504 784 508 785
rect 504 780 521 784
rect -431 715 335 719
rect -431 -66 -427 715
rect 418 714 515 718
rect -366 644 335 648
rect -366 -24 -362 644
rect 417 643 489 647
rect 327 604 331 608
rect 32 558 335 562
rect 417 557 423 561
rect 32 487 336 491
rect 418 486 422 490
rect 485 432 489 643
rect 511 608 515 714
rect 511 604 518 608
rect 515 568 516 572
rect 485 428 520 432
rect 32 416 335 420
rect 418 415 421 419
rect 32 345 335 349
rect 417 344 421 348
rect 1022 348 1031 352
rect 303 318 349 322
rect 133 277 193 281
rect 136 251 194 255
rect 136 248 140 251
rect 168 243 190 247
rect 168 181 172 243
rect 250 241 264 245
rect 303 230 307 318
rect 247 226 307 230
rect -7 178 1 180
rect -7 177 2 178
rect 137 177 142 181
rect 146 177 172 181
rect -7 176 1 177
rect 190 166 194 221
rect 121 162 194 166
rect 417 203 546 207
rect -7 105 5 109
rect 211 64 340 68
rect 140 35 141 39
rect 211 -24 215 64
rect 417 63 421 203
rect 430 194 546 198
rect -374 -28 215 -24
rect 233 -7 335 -3
rect 430 -4 434 194
rect -438 -67 -427 -66
rect 233 -67 237 -7
rect 418 -8 434 -4
rect 445 187 535 191
rect -438 -70 237 -67
rect -431 -71 237 -70
rect 309 -78 336 -74
rect 445 -75 449 187
rect 310 -100 314 -78
rect 418 -79 449 -75
rect 517 178 538 182
rect -500 -104 314 -100
rect -561 -149 335 -145
rect 517 -146 521 178
rect 1103 -126 1120 -122
rect -553 -1116 -549 -149
rect 417 -150 521 -146
rect -485 -1045 -481 -197
rect -429 -974 -425 -188
rect 326 -189 330 -185
rect -366 -903 -362 -191
rect 61 -235 335 -231
rect -267 -420 -262 -378
rect -267 -425 -255 -420
rect -260 -489 -255 -425
rect -204 -471 -201 -319
rect -149 -464 -145 -240
rect 57 -306 335 -302
rect 1110 -353 1126 -349
rect 56 -377 335 -373
rect 55 -448 335 -444
rect 948 -772 961 -768
rect -366 -907 352 -903
rect 430 -908 535 -904
rect -429 -978 349 -974
rect 431 -979 500 -975
rect -485 -1049 348 -1045
rect 431 -1050 479 -1046
rect -553 -1120 348 -1116
rect 430 -1121 459 -1117
rect 340 -1160 343 -1156
rect 76 -1206 348 -1202
rect 455 -1263 459 -1121
rect 475 -1192 479 -1050
rect 496 -1121 500 -979
rect 531 -1050 535 -908
rect 531 -1054 551 -1050
rect 618 -1055 628 -1051
rect 496 -1125 550 -1121
rect 619 -1126 631 -1122
rect 475 -1196 551 -1192
rect 619 -1197 629 -1193
rect 455 -1267 550 -1263
rect 618 -1268 627 -1264
rect 75 -1277 348 -1273
rect 77 -1348 348 -1344
rect 76 -1419 351 -1415
<< m2contact >>
rect 510 916 516 922
rect 511 744 516 749
rect 27 557 32 562
rect 423 557 428 562
rect 27 487 32 493
rect 422 486 427 491
rect 510 568 515 573
rect 26 415 32 421
rect 421 415 426 420
rect 510 390 515 395
rect 27 345 32 351
rect 421 344 426 349
rect 127 277 133 283
rect 546 203 551 208
rect 546 194 551 199
rect -366 -33 -361 -28
rect -431 -76 -425 -71
rect 535 186 540 191
rect -487 -109 -482 -104
rect 538 177 543 182
rect -429 -188 -424 -183
rect -487 -197 -481 -191
rect -367 -191 -361 -185
rect -149 -240 -144 -235
rect 55 -236 61 -230
rect 421 -237 426 -232
rect -206 -319 -201 -314
rect -268 -378 -262 -373
rect 51 -307 57 -301
rect 422 -309 428 -303
rect 50 -378 56 -372
rect 422 -380 428 -374
rect 49 -449 55 -443
rect 421 -451 427 -445
rect -149 -469 -143 -464
rect -206 -478 -200 -471
rect -261 -494 -255 -489
rect 69 -1208 76 -1200
rect 68 -1279 75 -1271
rect 70 -1350 77 -1342
rect 69 -1421 76 -1413
<< metal2 >>
rect 408 989 655 993
rect 127 901 344 905
rect 408 901 412 989
rect 1009 966 1028 970
rect 424 916 510 920
rect -309 560 27 561
rect -316 557 27 560
rect -487 -191 -483 -109
rect -429 -183 -425 -76
rect -366 -185 -362 -33
rect -316 -444 -312 557
rect -257 489 27 493
rect -257 -364 -253 489
rect -204 417 26 421
rect -204 -302 -200 417
rect -149 347 27 351
rect -149 -227 -145 347
rect 127 291 131 901
rect 424 562 428 916
rect 1024 790 1035 794
rect 434 744 511 748
rect 434 490 438 744
rect 1027 613 1040 617
rect 427 486 438 490
rect 451 568 510 572
rect 451 419 455 568
rect 1023 435 1036 439
rect 426 415 455 419
rect 473 390 510 394
rect 473 348 477 390
rect 426 344 477 348
rect 381 323 660 327
rect 540 187 555 190
rect 543 178 551 181
rect 338 146 343 152
rect 127 142 343 146
rect -161 -231 -145 -227
rect -149 -235 55 -231
rect -221 -306 51 -302
rect -206 -314 -202 -306
rect -272 -368 -253 -364
rect -257 -373 -253 -368
rect -262 -377 50 -373
rect -322 -448 49 -444
rect -316 -1415 -312 -448
rect -260 -1344 -256 -494
rect -205 -1273 -201 -478
rect -149 -1203 -145 -469
rect 291 -859 295 142
rect 339 108 343 142
rect 426 -236 517 -233
rect 428 -308 495 -305
rect 428 -379 468 -376
rect 427 -449 440 -446
rect 414 -708 418 -498
rect 437 -688 440 -449
rect 465 -676 468 -379
rect 492 -662 495 -308
rect 514 -648 517 -236
rect 514 -651 619 -648
rect 492 -665 616 -662
rect 465 -679 617 -676
rect 437 -691 619 -688
rect 414 -712 687 -708
rect 291 -863 358 -859
rect 419 -863 614 -859
rect 610 -1012 614 -863
rect -149 -1207 69 -1203
rect -205 -1277 68 -1273
rect -260 -1348 70 -1344
rect -316 -1419 69 -1415
<< m3contact >>
rect 338 152 343 157
rect 412 -498 418 -492
<< metal3 >>
rect 343 152 724 156
rect 133 -480 137 6
rect 133 -484 350 -480
rect 133 -1451 137 -484
rect 414 -492 418 -480
rect 616 -1451 620 -1299
rect 133 -1455 369 -1451
rect 425 -1455 620 -1451
use and_block  and_block_0
timestamp 1700077697
transform 1 0 560 0 1 -1093
box -18 -210 63 87
use enable_block  enable_block_2
timestamp 1700081456
transform 1 0 350 0 1 -1159
box -7 -296 85 300
use comp  comp_0
timestamp 1701515153
transform 1 0 905 0 1 -55
box -354 -732 209 261
use enable_block  enable_block_1
timestamp 1700081456
transform 1 0 337 0 1 -188
box -7 -296 85 300
use add_sub  add_sub_0
timestamp 1701536329
transform 1 0 671 0 1 841
box -156 -531 360 154
use enable_block  enable_block_0
timestamp 1700081456
transform 1 0 337 0 1 605
box -7 -296 85 300
use or  or_0
timestamp 1700071073
transform 1 0 184 0 1 217
box 1 0 70 65
use 2_4_decoder  2_4_decoder_0
timestamp 1700084785
transform 1 0 59 0 1 0
box -59 0 82 297
<< labels >>
rlabel metal1 -561 -149 -557 -145 3 a0
rlabel metal1 -500 -104 -496 -100 1 a1
rlabel metal1 -438 -70 -434 -66 1 a2
rlabel metal1 -374 -28 -370 -24 1 a3
rlabel metal2 -322 -448 -318 -444 1 b0
rlabel metal2 -272 -368 -268 -364 1 b1
rlabel metal2 -221 -306 -217 -302 1 b2
rlabel metal2 -161 -231 -157 -227 1 b3
rlabel metal1 623 -1268 627 -1264 1 ab3_and
rlabel metal1 625 -1197 629 -1193 1 ab2_and
rlabel metal1 627 -1126 631 -1122 1 ab1_and
rlabel metal1 624 -1055 628 -1051 1 ab0_and
rlabel metal1 957 -772 961 -768 1 a_eq_b
rlabel metal1 1122 -353 1126 -349 7 a_st_b
rlabel metal1 1116 -126 1120 -122 1 a_gt_b
rlabel metal2 1024 966 1028 970 1 sum1
rlabel metal2 1031 790 1035 794 1 sum2
rlabel metal2 1036 613 1040 617 1 sum3
rlabel metal2 1032 435 1036 439 1 sum4
rlabel metal1 1027 348 1031 352 1 carry
rlabel metal1 -7 176 -3 180 1 s1
rlabel metal1 -7 105 -3 109 1 s0
rlabel metal2 408 989 412 993 5 vdd
rlabel metal2 449 323 453 327 1 gnd
rlabel metal1 148 251 151 255 1 check1
rlabel metal1 159 177 162 181 1 check2
rlabel polysilicon 149 107 151 109 1 check3
rlabel polysilicon 142 -8 144 -6 1 check4
<< end >>
