magic
tech scmos
timestamp 1700071073
<< metal1 >>
rect 5 60 6 64
rect 6 34 7 38
rect 6 26 7 30
rect 34 25 45 29
rect 69 24 70 28
rect 6 0 7 4
<< m2contact >>
rect 23 60 28 65
rect 44 47 49 52
rect 44 8 49 13
rect 24 0 29 5
<< metal2 >>
rect 28 60 48 64
rect 44 52 48 60
rect 44 4 48 8
rect 29 0 48 4
use inverter  inverter_0
timestamp 1700050252
transform 1 0 76 0 1 43
box -32 -34 -7 8
use nor  nor_0
timestamp 1700050543
transform 1 0 1 0 1 40
box 0 -40 37 24
<< end >>
