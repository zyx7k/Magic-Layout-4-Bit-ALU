magic
tech scmos
timestamp 1700050467
<< nwell >>
rect 0 0 52 18
<< ntransistor >>
rect 12 -37 14 -31
rect 22 -37 24 -31
rect 30 -37 32 -31
rect 38 -37 40 -31
<< ptransistor >>
rect 12 6 14 12
rect 22 6 24 12
rect 30 6 32 12
rect 38 6 40 12
<< ndiffusion >>
rect 6 -32 12 -31
rect 6 -37 7 -32
rect 11 -37 12 -32
rect 14 -37 22 -31
rect 24 -37 30 -31
rect 32 -37 38 -31
rect 40 -36 43 -31
rect 47 -36 48 -31
rect 40 -37 48 -36
<< pdiffusion >>
rect 6 7 7 12
rect 11 7 12 12
rect 6 6 12 7
rect 14 11 22 12
rect 14 6 17 11
rect 21 6 22 11
rect 24 7 25 12
rect 29 7 30 12
rect 24 6 30 7
rect 32 11 38 12
rect 32 6 33 11
rect 37 6 38 11
rect 40 7 41 12
rect 45 7 46 12
rect 40 6 46 7
<< ndcontact >>
rect 7 -37 11 -32
rect 43 -36 47 -31
<< pdcontact >>
rect 7 7 11 12
rect 17 6 21 11
rect 25 7 29 12
rect 33 6 37 11
rect 41 7 45 12
<< polysilicon >>
rect 12 12 14 15
rect 22 12 24 15
rect 30 12 32 15
rect 38 12 40 15
rect 12 -2 14 6
rect 12 -31 14 -6
rect 22 -10 24 6
rect 22 -31 24 -14
rect 30 -17 32 6
rect 30 -31 32 -21
rect 38 -24 40 6
rect 38 -31 40 -28
rect 12 -40 14 -37
rect 22 -40 24 -37
rect 30 -40 32 -37
rect 38 -40 40 -37
<< polycontact >>
rect 10 -6 14 -2
rect 20 -14 24 -10
rect 28 -21 32 -17
rect 36 -28 40 -24
<< metal1 >>
rect 0 20 52 24
rect 7 12 11 20
rect 25 12 29 20
rect 41 12 45 20
rect 17 -2 21 6
rect 33 -2 37 6
rect 6 -6 10 -2
rect 17 -6 47 -2
rect 6 -14 20 -10
rect 6 -21 28 -17
rect 6 -28 36 -24
rect 43 -31 47 -6
rect 7 -42 11 -37
rect 6 -46 48 -42
<< end >>
