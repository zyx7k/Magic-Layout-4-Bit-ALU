magic
tech scmos
timestamp 1701515153
<< polysilicon >>
rect -179 214 29 216
rect -235 172 -233 181
rect -235 170 -207 172
rect -179 135 -177 214
rect -204 133 -177 135
rect -174 209 -11 211
rect 27 210 29 214
rect -269 126 -216 128
rect -280 6 -278 20
rect -269 4 -267 126
rect -174 100 -172 209
rect -204 98 -172 100
rect -169 204 -27 206
rect -257 90 -215 92
rect -257 -6 -255 90
rect -169 65 -167 204
rect -204 63 -167 65
rect -164 199 -88 201
rect -248 56 -215 58
rect -248 -6 -246 56
rect -164 29 -162 199
rect -204 27 -162 29
rect -166 11 -123 13
rect -150 3 -144 5
rect -150 2 -148 3
rect -125 3 -123 11
rect -166 0 -148 2
rect -90 -129 -88 199
rect -29 6 -27 204
rect -13 104 -11 209
rect -6 110 -4 199
rect 29 122 100 124
rect -6 108 11 110
rect -13 102 22 104
rect -4 95 7 97
rect 30 18 95 20
rect -19 11 39 13
rect -29 4 31 6
rect -36 -93 -34 3
rect -5 -4 24 -2
rect -21 -14 17 -12
rect 93 -42 95 18
rect 98 -35 100 122
rect 98 -38 109 -35
rect 93 -46 98 -42
rect 90 -52 109 -50
rect 90 -86 92 -52
rect 18 -88 92 -86
rect -36 -95 43 -93
rect -5 -104 36 -102
rect -5 -113 29 -111
rect -5 -122 22 -120
rect -90 -131 15 -129
rect -280 -170 -278 -158
rect -269 -170 -267 -158
rect -257 -171 -255 -158
rect -248 -181 -246 -158
rect -166 -166 -122 -164
rect -151 -173 -144 -171
rect -166 -175 -149 -173
rect -124 -172 -122 -166
rect -100 -166 -78 -164
rect 96 -215 98 -56
rect 22 -217 98 -215
rect -57 -225 26 -223
rect -334 -432 -332 -328
rect -326 -394 -324 -328
rect -280 -350 -278 -329
rect -269 -350 -267 -329
rect -257 -350 -255 -329
rect -248 -346 -246 -329
rect -164 -341 -123 -339
rect -125 -346 -123 -341
rect -115 -341 -71 -339
rect -164 -348 -133 -346
rect -204 -389 -164 -387
rect -326 -396 -216 -394
rect -204 -428 -170 -426
rect -334 -434 -216 -432
rect -204 -466 -176 -464
rect -346 -474 -216 -472
rect -207 -628 -205 -503
rect -178 -614 -176 -466
rect -172 -600 -170 -428
rect -166 -586 -164 -389
rect -75 -435 -65 -433
rect -118 -532 -116 -521
rect -118 -534 -65 -532
rect -57 -586 -55 -225
rect -166 -588 -55 -586
rect -52 -233 18 -231
rect -52 -594 -50 -233
rect 68 -265 112 -263
rect 68 -296 70 -265
rect 29 -298 70 -296
rect 75 -273 102 -271
rect -103 -596 -50 -594
rect -47 -305 28 -303
rect -47 -600 -45 -305
rect -172 -602 -45 -600
rect -42 -313 21 -311
rect -42 -608 -40 -313
rect -7 -322 14 -320
rect 75 -401 77 -273
rect 29 -403 77 -401
rect 83 -279 93 -277
rect -103 -610 -40 -608
rect -37 -410 39 -408
rect -37 -614 -35 -410
rect -178 -616 -35 -614
rect -32 -418 31 -416
rect -32 -622 -30 -418
rect -5 -427 24 -425
rect -5 -435 17 -433
rect 83 -513 85 -279
rect 18 -515 85 -513
rect 99 -287 112 -285
rect -7 -522 43 -520
rect -7 -530 36 -528
rect -103 -624 -30 -622
rect -27 -538 29 -536
rect -27 -628 -25 -538
rect -207 -630 -25 -628
rect -22 -547 22 -545
rect -22 -633 -20 -547
rect -6 -554 15 -552
rect -98 -635 -20 -633
rect -98 -636 -96 -635
rect -103 -638 -96 -636
rect 99 -641 101 -287
rect 22 -643 101 -641
<< polycontact >>
rect -236 181 -232 185
rect -207 169 -203 173
rect -208 132 -204 136
rect -281 20 -277 24
rect -281 2 -277 6
rect -216 125 -212 129
rect -208 97 -204 101
rect -270 0 -266 4
rect -215 89 -211 93
rect -208 63 -204 67
rect -215 55 -211 59
rect -208 26 -204 30
rect -170 11 -166 15
rect -170 0 -166 4
rect -144 2 -140 6
rect -125 -1 -121 3
rect -258 -10 -254 -6
rect -249 -10 -245 -6
rect -38 3 -34 7
rect 26 206 30 210
rect -7 199 -3 203
rect 25 121 29 125
rect 11 108 15 112
rect 22 100 26 104
rect -8 94 -4 98
rect 7 94 11 98
rect 26 17 30 21
rect -23 11 -19 15
rect 39 10 43 14
rect 31 3 35 7
rect -9 -5 -5 -1
rect 24 -5 28 -1
rect -25 -16 -21 -12
rect 17 -16 21 -12
rect 109 -39 113 -35
rect 98 -46 102 -42
rect 14 -89 18 -85
rect 109 -53 113 -49
rect 43 -96 47 -92
rect -9 -106 -5 -102
rect 36 -105 40 -101
rect -9 -115 -5 -111
rect 29 -114 33 -110
rect -9 -124 -5 -120
rect 22 -123 26 -119
rect 15 -132 19 -128
rect -281 -158 -277 -154
rect -270 -158 -266 -154
rect -258 -158 -254 -154
rect -249 -158 -245 -154
rect -281 -174 -277 -170
rect -270 -174 -266 -170
rect -258 -175 -254 -171
rect -170 -166 -166 -162
rect -170 -175 -166 -171
rect -144 -174 -140 -170
rect -104 -167 -100 -163
rect -78 -167 -74 -163
rect -125 -176 -121 -172
rect -249 -185 -245 -181
rect 18 -218 22 -214
rect 98 -60 102 -56
rect -335 -328 -331 -324
rect -327 -328 -323 -324
rect -281 -329 -277 -325
rect -270 -329 -266 -325
rect -258 -329 -254 -325
rect -249 -329 -245 -325
rect -168 -341 -164 -337
rect -119 -342 -115 -338
rect -71 -341 -67 -337
rect -249 -350 -245 -346
rect -168 -350 -164 -346
rect -133 -350 -129 -346
rect -125 -350 -121 -346
rect -281 -354 -277 -350
rect -270 -354 -266 -350
rect -258 -354 -254 -350
rect -208 -390 -204 -386
rect -216 -397 -212 -393
rect -208 -429 -204 -425
rect -216 -435 -212 -431
rect -208 -467 -204 -463
rect -350 -474 -346 -470
rect -216 -475 -212 -471
rect -208 -503 -204 -499
rect -79 -437 -75 -433
rect -65 -437 -61 -433
rect -119 -521 -115 -517
rect -65 -535 -61 -531
rect 26 -226 30 -222
rect -107 -596 -103 -592
rect 18 -235 22 -231
rect 25 -299 29 -295
rect 112 -266 116 -262
rect 102 -273 106 -269
rect 28 -307 32 -303
rect -107 -610 -103 -606
rect 21 -315 25 -311
rect -11 -322 -7 -318
rect 14 -324 18 -320
rect 25 -404 29 -400
rect 39 -411 43 -407
rect -107 -624 -103 -620
rect 31 -419 35 -415
rect -9 -429 -5 -425
rect 24 -428 28 -424
rect -9 -437 -5 -433
rect 17 -437 21 -433
rect 14 -516 18 -512
rect 93 -281 97 -277
rect 112 -287 116 -283
rect -11 -522 -7 -518
rect 43 -523 47 -519
rect -11 -530 -7 -526
rect 36 -531 40 -527
rect 29 -539 33 -535
rect 22 -548 26 -544
rect -10 -556 -6 -552
rect 15 -556 19 -552
rect -107 -638 -103 -634
rect 18 -644 22 -640
<< metal1 >>
rect -350 -338 -347 231
rect -342 227 -339 256
rect -335 -162 -331 240
rect -327 227 -324 249
rect -295 15 -291 249
rect -232 197 -228 256
rect -232 193 -121 197
rect -281 185 -128 189
rect -281 24 -277 185
rect -161 171 -157 177
rect -133 174 -128 185
rect -125 177 -121 193
rect -207 160 -203 169
rect -207 158 -204 160
rect -223 118 -219 138
rect -208 136 -204 138
rect -212 125 -203 129
rect -185 122 -181 139
rect -223 82 -219 105
rect -208 101 -204 103
rect -211 89 -203 93
rect -185 84 -181 104
rect -223 47 -219 65
rect -211 55 -203 59
rect -185 48 -181 67
rect -161 51 -157 56
rect -96 30 -92 62
rect -295 11 -170 15
rect -119 13 -115 17
rect -281 -154 -277 2
rect -266 0 -170 4
rect -270 -154 -266 0
rect -161 -2 -157 4
rect -140 3 -128 6
rect -140 2 -130 3
rect -96 -4 -92 23
rect -37 7 -34 233
rect -23 15 -20 233
rect -7 203 -3 233
rect -1 186 3 187
rect 18 182 22 233
rect 26 181 30 206
rect 61 185 65 191
rect 15 108 33 112
rect -12 95 -8 98
rect 11 94 19 98
rect 15 90 19 94
rect 22 89 26 100
rect 29 91 33 108
rect -12 -4 -9 -1
rect -258 -154 -254 -10
rect -249 -154 -245 -10
rect -78 -15 -25 -12
rect -78 -111 -75 -15
rect -1 -14 3 -13
rect 24 -14 28 -5
rect 31 -14 35 3
rect 39 -14 43 10
rect 65 -12 112 -8
rect 102 -46 113 -42
rect 102 -60 113 -56
rect 190 -71 204 -67
rect -16 -105 -9 -102
rect -161 -124 -157 -120
rect -96 -136 -92 -112
rect -78 -114 -9 -111
rect -118 -139 -114 -136
rect -335 -166 -170 -162
rect -119 -163 -115 -159
rect -335 -324 -331 -166
rect -119 -167 -104 -163
rect -327 -324 -323 -320
rect -281 -325 -277 -174
rect -270 -325 -266 -174
rect -254 -175 -170 -171
rect -258 -325 -254 -175
rect -161 -177 -157 -172
rect -140 -173 -128 -170
rect -140 -174 -132 -173
rect -96 -182 -92 -156
rect -78 -163 -75 -114
rect -71 -123 -9 -120
rect -249 -325 -245 -185
rect -161 -299 -157 -295
rect -96 -311 -92 -291
rect -350 -341 -168 -338
rect -119 -338 -115 -334
rect -350 -470 -347 -341
rect -245 -349 -168 -346
rect -281 -591 -277 -354
rect -270 -605 -266 -354
rect -258 -619 -254 -354
rect -249 -631 -246 -350
rect -133 -353 -128 -350
rect -125 -353 -121 -350
rect -211 -358 -203 -354
rect -161 -358 -157 -354
rect -96 -358 -92 -330
rect -207 -359 -203 -358
rect -223 -400 -219 -380
rect -208 -386 -204 -384
rect -212 -397 -203 -393
rect -207 -398 -203 -397
rect -185 -398 -181 -379
rect -223 -435 -219 -419
rect -208 -425 -204 -423
rect -212 -435 -203 -432
rect -185 -435 -181 -418
rect -78 -433 -75 -167
rect -207 -438 -204 -435
rect -223 -477 -219 -456
rect -208 -463 -204 -460
rect -212 -474 -203 -471
rect -212 -475 -205 -474
rect -185 -477 -181 -455
rect -161 -490 -157 -475
rect -96 -490 -92 -472
rect -161 -494 -134 -490
rect -208 -499 -204 -498
rect -119 -517 -115 -514
rect -78 -523 -75 -437
rect -71 -337 -68 -123
rect -1 -134 3 -85
rect 59 -86 119 -82
rect 15 -138 19 -132
rect 22 -138 26 -123
rect 29 -138 33 -114
rect 36 -138 40 -105
rect 43 -138 47 -96
rect 18 -214 22 -213
rect 26 -239 30 -226
rect 107 -236 110 -235
rect 61 -240 110 -236
rect 106 -273 116 -269
rect 101 -277 116 -276
rect 97 -280 116 -277
rect 97 -281 101 -280
rect 193 -298 209 -294
rect -17 -322 -11 -319
rect 14 -334 18 -324
rect 21 -334 25 -315
rect 28 -335 32 -307
rect 51 -313 121 -309
rect -71 -519 -68 -341
rect -13 -428 -9 -425
rect -61 -436 -9 -433
rect 17 -446 21 -437
rect 24 -446 28 -428
rect 31 -446 35 -419
rect 39 -446 43 -411
rect -71 -522 -11 -519
rect -229 -596 -107 -593
rect -229 -610 -107 -607
rect -229 -624 -107 -621
rect -229 -636 -107 -633
rect -110 -637 -107 -636
rect -86 -710 -83 -644
rect -78 -703 -75 -528
rect -71 -696 -68 -522
rect -15 -530 -11 -527
rect -65 -688 -62 -535
rect -13 -555 -10 -552
rect -1 -565 3 -508
rect 15 -565 19 -556
rect 22 -565 26 -548
rect 29 -565 33 -539
rect 36 -565 40 -531
rect 43 -565 47 -523
rect -65 -689 -51 -688
rect -65 -692 -52 -689
rect -71 -700 -52 -696
rect -78 -706 -50 -703
rect -78 -707 -51 -706
rect -86 -712 -50 -710
rect -86 -714 -52 -712
rect 16 -717 48 -713
rect 15 -732 25 -728
<< m2contact >>
rect -344 256 -339 261
rect -233 256 -228 261
rect -352 231 -347 236
rect -327 249 -322 254
rect -296 249 -291 254
rect -336 240 -331 245
rect -343 222 -338 227
rect -328 222 -323 227
rect -37 233 -32 238
rect -23 233 -18 238
rect -7 233 -2 238
rect 18 233 23 238
rect -161 177 -156 182
rect -97 173 -92 178
rect -223 161 -218 166
rect -185 161 -180 166
rect -161 46 -156 51
rect -119 41 -114 46
rect -135 36 -130 41
rect -161 4 -156 9
rect -119 7 -113 13
rect -1 187 4 192
rect 61 191 66 196
rect -17 95 -12 100
rect -1 87 4 92
rect 61 96 66 101
rect -17 -6 -12 -1
rect -1 -13 4 -8
rect 64 -8 69 -3
rect -2 -85 3 -80
rect -21 -107 -16 -102
rect -161 -129 -156 -124
rect -135 -140 -130 -135
rect -119 -136 -114 -131
rect -328 -320 -323 -315
rect -161 -172 -156 -167
rect -161 -304 -156 -299
rect -119 -310 -114 -305
rect -135 -315 -130 -310
rect -282 -596 -277 -591
rect -271 -610 -266 -605
rect -259 -624 -254 -619
rect -216 -358 -211 -353
rect -161 -354 -156 -349
rect -119 -490 -114 -485
rect -223 -504 -218 -499
rect -186 -503 -181 -498
rect -135 -520 -130 -515
rect -97 -519 -92 -514
rect 54 -86 59 -81
rect 68 -128 73 -123
rect -22 -322 -17 -317
rect -3 -330 3 -325
rect 45 -314 51 -308
rect 61 -325 66 -320
rect -18 -430 -13 -425
rect -2 -442 3 -437
rect 65 -436 70 -431
rect -79 -528 -74 -523
rect -234 -596 -229 -591
rect -234 -610 -229 -605
rect -234 -624 -229 -619
rect -251 -636 -246 -631
rect -234 -636 -229 -631
rect -86 -644 -81 -639
rect -20 -530 -15 -525
rect -18 -557 -13 -552
rect 68 -555 73 -550
rect 2 -644 7 -639
rect 25 -732 30 -727
<< metal2 >>
rect -354 258 -344 261
rect -339 258 -233 261
rect -228 258 21 261
rect -354 249 -327 252
rect -322 249 -296 252
rect -291 249 -4 252
rect -354 242 -336 245
rect -331 242 -20 245
rect -23 238 -20 242
rect -7 238 -4 249
rect 18 238 21 258
rect -354 233 -352 236
rect -347 233 -37 236
rect -223 225 73 229
rect -342 -355 -339 222
rect -327 -315 -324 222
rect -223 166 -219 225
rect -161 182 -157 225
rect -1 192 3 225
rect 61 196 65 201
rect -96 178 -92 182
rect -185 166 -181 170
rect -86 95 -17 98
rect -119 46 -115 47
rect -161 41 -157 46
rect -161 37 -135 41
rect -161 9 -157 37
rect -86 10 -83 95
rect -1 92 3 150
rect 61 101 65 150
rect -113 7 -83 10
rect -86 -1 -83 7
rect -86 -4 -17 -1
rect -86 -102 -83 -4
rect 0 -8 4 46
rect 62 41 69 45
rect 65 -3 69 41
rect 64 -70 72 -66
rect 3 -85 54 -81
rect -86 -105 -21 -102
rect -161 -136 -157 -129
rect -119 -131 -115 -127
rect -161 -140 -135 -136
rect -161 -167 -157 -140
rect -161 -310 -157 -304
rect -119 -305 -115 -303
rect -161 -314 -135 -310
rect -161 -349 -157 -314
rect -86 -319 -83 -105
rect 68 -123 72 -70
rect -1 -308 3 -271
rect -1 -312 45 -308
rect -86 -322 -22 -319
rect -342 -358 -216 -355
rect -86 -425 -83 -322
rect -1 -325 3 -312
rect 61 -320 65 -271
rect -86 -428 -18 -425
rect -119 -485 -115 -484
rect -292 -596 -282 -593
rect -277 -596 -234 -593
rect -292 -610 -271 -607
rect -266 -610 -234 -607
rect -292 -624 -259 -621
rect -254 -624 -234 -621
rect -292 -636 -251 -633
rect -246 -636 -234 -633
rect -223 -653 -219 -504
rect -185 -508 -181 -503
rect -134 -653 -130 -520
rect -96 -524 -92 -519
rect -86 -552 -83 -428
rect -1 -437 3 -375
rect 61 -380 69 -376
rect 65 -431 69 -380
rect 65 -498 72 -494
rect -74 -528 -20 -525
rect 68 -550 72 -498
rect -86 -555 -18 -552
rect -86 -639 -83 -555
rect 3 -653 7 -644
rect -223 -657 30 -653
rect 26 -727 30 -657
<< m3contact >>
rect 61 201 66 206
rect -97 182 -92 187
rect -185 170 -180 175
rect -186 -513 -181 -508
rect -97 -529 -92 -524
rect 65 -629 72 -622
rect 0 -666 5 -661
<< metal3 >>
rect -185 219 73 223
rect -185 175 -181 219
rect -96 187 -92 219
rect 61 206 65 219
rect -185 -648 -181 -513
rect -95 -648 -92 -529
rect 67 -648 72 -629
rect -185 -651 72 -648
rect 0 -661 3 -651
use and4  and4_2
timestamp 1700071032
transform 1 0 -52 0 1 -728
box -6 -4 72 67
use and5  and5_1
timestamp 1700071052
transform 0 1 -1 -1 0 -556
box -1 0 86 74
use inverter  inverter_3
timestamp 1700050252
transform 0 1 -100 -1 0 -522
box -32 -34 -7 8
use xor  xor_3
timestamp 1700050706
transform 0 1 -129 -1 0 -371
box -18 -32 113 37
use inverter  inverter_4
timestamp 1700050252
transform 0 1 -189 -1 0 -506
box -32 -34 -7 8
use and4  and4_1
timestamp 1700071032
transform 0 1 3 -1 0 -442
box -6 -4 72 67
use inverter  inverter_7
timestamp 1700050252
transform 0 1 -189 -1 0 -391
box -32 -34 -7 8
use inverter  inverter_6
timestamp 1700050252
transform 0 1 -189 -1 0 -430
box -32 -34 -7 8
use inverter  inverter_5
timestamp 1700050252
transform 0 1 -189 -1 0 -467
box -32 -34 -7 8
use and3  and3_1
timestamp 1700071010
transform 0 1 -1 -1 0 -325
box 0 -1 77 67
use inverter  inverter_2
timestamp 1700050252
transform 0 1 -100 -1 0 -342
box -32 -34 -7 8
use xor  xor_2
timestamp 1700050706
transform 0 1 -129 -1 0 -190
box -18 -32 113 37
use and  and_1
timestamp 1700070968
transform 0 1 -1 -1 0 -230
box 0 0 67 67
use and5  and5_0
timestamp 1700071052
transform 0 1 -1 -1 0 -129
box -1 0 86 74
use or4  or4_1
timestamp 1700071115
transform 1 0 112 0 1 -313
box -2 0 85 78
use inverter  inverter_1
timestamp 1700050252
transform 0 1 -100 -1 0 -168
box -32 -34 -7 8
use xor  xor_1
timestamp 1700050706
transform 0 1 -129 -1 0 -15
box -18 -32 113 37
use and4  and4_0
timestamp 1700071032
transform 0 1 3 -1 0 -14
box -6 -4 72 67
use or4  or4_0
timestamp 1700071115
transform 1 0 109 0 1 -86
box -2 0 85 78
use inverter  inverter_0
timestamp 1700050252
transform 0 1 -100 -1 0 9
box -32 -34 -7 8
use inverter  inverter_11
timestamp 1700050252
transform 0 1 -189 -1 0 23
box -32 -34 -7 8
use xor  xor_0
timestamp 1700050706
transform 0 1 -129 -1 0 160
box -18 -32 113 37
use and3  and3_0
timestamp 1700071010
transform 0 1 0 -1 0 96
box 0 -1 77 67
use inverter  inverter_10
timestamp 1700050252
transform 0 1 -189 -1 0 58
box -32 -34 -7 8
use inverter  inverter_9
timestamp 1700050252
transform 0 1 -189 -1 0 94
box -32 -34 -7 8
use inverter  inverter_8
timestamp 1700050252
transform 0 1 -189 -1 0 129
box -32 -34 -7 8
use and  and_0
timestamp 1700070968
transform 0 1 -1 -1 0 191
box 0 0 67 67
<< end >>
