magic
tech scmos
timestamp 1699993993
<< nwell >>
rect 0 0 49 17
<< ntransistor >>
rect 11 -28 13 -23
rect 19 -28 21 -23
rect 27 -28 29 -23
<< ptransistor >>
rect 11 6 13 11
rect 19 6 21 11
rect 27 6 29 11
<< ndiffusion >>
rect 10 -28 11 -23
rect 13 -28 14 -23
rect 18 -28 19 -23
rect 21 -28 22 -23
rect 26 -28 27 -23
rect 29 -28 33 -23
<< pdiffusion >>
rect 10 6 11 11
rect 13 6 19 11
rect 21 6 27 11
rect 29 6 33 11
<< ndcontact >>
rect 6 -28 10 -23
rect 14 -28 18 -23
rect 22 -28 26 -23
rect 33 -28 37 -23
<< pdcontact >>
rect 6 6 10 11
rect 33 6 37 11
<< polysilicon >>
rect 11 11 13 14
rect 19 11 21 14
rect 27 11 29 14
rect 11 -23 13 6
rect 19 -8 21 6
rect 27 -1 29 6
rect 19 -23 21 -12
rect 27 -23 29 -5
rect 11 -31 13 -28
rect 19 -31 21 -28
rect 27 -31 29 -28
<< polycontact >>
rect 7 -19 11 -15
rect 26 -5 30 -1
rect 18 -12 22 -8
<< metal1 >>
rect 0 18 49 22
rect 6 11 10 18
rect 0 -5 26 -1
rect 0 -12 18 -8
rect 33 -15 37 6
rect 0 -19 7 -15
rect 14 -19 37 -15
rect 14 -23 18 -19
rect 33 -23 37 -19
rect 6 -32 10 -28
rect 22 -32 26 -28
rect 0 -36 48 -32
<< labels >>
rlabel metal1 4 -18 6 -16 3 a
rlabel metal1 4 -11 6 -9 3 b
rlabel metal1 4 -4 6 -2 3 c
rlabel metal1 7 -32 9 -30 1 gnd
rlabel metal1 7 18 9 20 5 vdd
rlabel metal1 34 -18 36 -16 1 out
<< end >>
