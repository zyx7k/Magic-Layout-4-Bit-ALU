magic
tech scmos
timestamp 1700050393
<< nwell >>
rect -8 -3 37 14
<< ntransistor >>
rect 5 -38 7 -33
rect 13 -38 15 -33
rect 21 -38 23 -33
<< ptransistor >>
rect 5 3 7 8
rect 13 3 15 8
rect 21 3 23 8
<< ndiffusion >>
rect -2 -34 5 -33
rect -2 -38 -1 -34
rect 3 -38 5 -34
rect 7 -38 13 -33
rect 15 -38 21 -33
rect 23 -37 26 -33
rect 30 -37 31 -33
rect 23 -38 31 -37
<< pdiffusion >>
rect -2 4 -1 8
rect 3 4 5 8
rect -2 3 5 4
rect 7 7 13 8
rect 7 3 8 7
rect 12 3 13 7
rect 15 4 16 8
rect 20 4 21 8
rect 15 3 21 4
rect 23 7 31 8
rect 23 3 26 7
rect 30 3 31 7
<< ndcontact >>
rect -1 -38 3 -34
rect 26 -37 30 -33
<< pdcontact >>
rect -1 4 3 8
rect 8 3 12 7
rect 16 4 20 8
rect 26 3 30 7
<< polysilicon >>
rect 5 8 7 12
rect 13 8 15 12
rect 21 8 23 12
rect 5 -27 7 3
rect 13 -20 15 3
rect 21 -13 23 3
rect 5 -33 7 -31
rect 13 -33 15 -24
rect 21 -33 23 -17
rect 5 -41 7 -38
rect 13 -41 15 -38
rect 21 -41 23 -38
<< polycontact >>
rect 19 -17 23 -13
rect 11 -24 15 -20
rect 3 -31 7 -27
<< metal1 >>
rect -7 16 33 20
rect -1 8 3 16
rect 16 8 20 16
rect 8 -5 12 3
rect 26 -5 30 3
rect 8 -9 30 -5
rect -2 -17 19 -13
rect 26 -15 30 -9
rect 26 -19 33 -15
rect -2 -24 11 -20
rect -2 -31 3 -27
rect 26 -33 30 -19
rect -1 -42 3 -38
rect -2 -46 22 -42
<< end >>
