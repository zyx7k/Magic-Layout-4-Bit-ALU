magic
tech scmos
timestamp 1700050600
<< nwell >>
rect 0 0 60 18
<< ntransistor >>
rect 14 -44 16 -39
rect 23 -44 25 -39
rect 33 -44 35 -39
rect 43 -44 45 -39
<< ptransistor >>
rect 14 6 16 12
rect 23 6 25 12
rect 33 6 35 12
rect 43 6 45 12
<< ndiffusion >>
rect 7 -40 14 -39
rect 7 -44 8 -40
rect 12 -44 14 -40
rect 16 -40 23 -39
rect 16 -44 18 -40
rect 22 -44 23 -40
rect 25 -40 33 -39
rect 25 -44 27 -40
rect 31 -44 33 -40
rect 35 -40 43 -39
rect 35 -44 38 -40
rect 42 -44 43 -40
rect 45 -40 51 -39
rect 45 -44 46 -40
rect 50 -44 51 -40
<< pdiffusion >>
rect 6 7 7 12
rect 11 7 14 12
rect 6 6 14 7
rect 16 6 23 12
rect 25 6 33 12
rect 35 6 43 12
rect 45 11 54 12
rect 45 6 49 11
rect 53 6 54 11
<< ndcontact >>
rect 8 -44 12 -40
rect 18 -44 22 -40
rect 27 -44 31 -40
rect 38 -44 42 -40
rect 46 -44 50 -40
<< pdcontact >>
rect 7 7 11 12
rect 49 6 53 11
<< polysilicon >>
rect 14 12 16 15
rect 23 12 25 15
rect 33 12 35 15
rect 43 12 45 15
rect 14 -16 16 6
rect 23 -9 25 6
rect 33 -2 35 6
rect 14 -39 16 -20
rect 23 -39 25 -13
rect 33 -39 35 -6
rect 43 -23 45 6
rect 43 -39 45 -27
rect 14 -47 16 -44
rect 23 -47 25 -44
rect 33 -47 35 -44
rect 43 -47 45 -44
<< polycontact >>
rect 31 -6 35 -2
rect 22 -13 26 -9
rect 12 -20 16 -16
rect 42 -27 46 -23
<< metal1 >>
rect 0 21 60 25
rect 7 12 11 21
rect 7 -6 31 -2
rect 7 -13 22 -9
rect 49 -15 53 6
rect 7 -20 12 -16
rect 49 -19 55 -15
rect 7 -27 42 -23
rect 49 -32 53 -19
rect 18 -36 53 -32
rect 18 -40 22 -36
rect 38 -40 42 -36
rect 8 -49 12 -44
rect 27 -49 31 -44
rect 46 -49 50 -44
rect 7 -53 51 -49
<< end >>
