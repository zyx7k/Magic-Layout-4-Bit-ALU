magic
tech scmos
timestamp 1700050252
<< nwell >>
rect -32 -12 -8 4
<< ntransistor >>
rect -21 -26 -19 -22
<< ptransistor >>
rect -21 -6 -19 -2
<< ndiffusion >>
rect -22 -26 -21 -22
rect -19 -26 -18 -22
<< pdiffusion >>
rect -22 -6 -21 -2
rect -19 -6 -18 -2
<< ndcontact >>
rect -26 -26 -22 -22
rect -18 -26 -14 -22
<< pdcontact >>
rect -26 -6 -22 -2
rect -18 -6 -14 -2
<< polysilicon >>
rect -21 -2 -19 1
rect -21 -15 -19 -6
rect -25 -17 -19 -15
rect -21 -22 -19 -17
rect -21 -29 -19 -26
<< polycontact >>
rect -29 -18 -25 -14
<< metal1 >>
rect -32 4 -8 8
rect -26 -2 -22 4
rect -32 -18 -29 -14
rect -18 -15 -14 -6
rect -18 -19 -7 -15
rect -18 -22 -14 -19
rect -26 -30 -22 -26
rect -32 -34 -7 -30
<< end >>
