magic
tech scmos
timestamp 1700071115
<< metal1 >>
rect -2 74 0 78
rect 4 47 7 51
rect 4 40 7 44
rect 4 33 7 37
rect 4 26 7 30
rect 50 18 58 20
rect 49 16 58 18
rect 83 15 85 19
rect 5 0 7 4
rect 50 0 59 4
<< m2contact >>
rect 55 73 60 78
rect 64 38 69 43
<< metal2 >>
rect 60 74 68 78
rect 64 43 68 74
use inverter  inverter_0
timestamp 1700050252
transform 1 0 90 0 1 34
box -32 -34 -7 8
use nor4  nor4_0
timestamp 1700050600
transform 1 0 0 0 1 53
box 0 -53 60 25
<< end >>
